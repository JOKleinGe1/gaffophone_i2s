module i2s(
endmodule

